library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;



entity alpha_computation_even is 
	
	generic(
		W_bits			: positive := 32; -- size of word
		F_bits			: positive := 16); -- number of newton's iterations
		
	port(	clock		: in std_logic;
		beta_even	: in unsigned(W_bits-1 downto 0);
		alpha_even	: out unsigned(W_bits-1 downto 0));
		
end entity alpha_computation_even;
 	


architecture alpha_even_comp_arch of alpha_computation_even is

	-- Beta Even Alpha = -2*B + .5*B

	signal beta_one		: unsigned(W_bits-1 downto 0);
	signal beta_two		: unsigned(W_bits-1 downto 0);
	begin
	

	process(clock)

	begin
		if(rising_edge(clock)) then
		
		beta_one <= beta_even;
		beta_two <= beta_even;

		beta_one <= shift_left(beta_even,1);

		beta_two <= shift_right(beta_even,1);
		
		alpha_even <= beta_two - beta_one;
		
		end if;

	end process;
	
end architecture;
