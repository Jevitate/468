library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity rsqrt is 
	
	generic(
		W_bits			: positive := 32; -- size of word
		F_bits			: positive := 16; -- number of fractional bits
		N_iterations		: positive := 3); -- number of newton's iterations
		
	port(	clock	: in std_logic;
		x	: in std_logic_vector(W_bits-1 downto 0);
		x_test	: out std_logic_vector(W_bits-1 downto 0);
		y_test	: out std_logic_vector(W_bits-1 downto 0);
		y_0	: in std_logic_vector(W_bits-1 downto 0);
		y	: out std_logic_vector(W_bits-1 downto 0));
		
end entity rsqrt;

--0000 0000 0000 0000 . 0000 0000 0000 0000

architecture rsqrt_arch of rsqrt is

	signal arithimetric 		: unsigned(W_bits-1 downto 0);
	signal three			: unsigned(W_bits-1 downto 0); -- W - F - 00s, 2 1s,

	signal yn_squared		: unsigned(2*W_bits-1 downto 0);
	signal yn_squared_resized	: unsigned(W_bits-1 downto 0);

	signal x_yn_2			: unsigned(2*W_bits-1 downto 0);
	signal x_yn_2_resized		: unsigned(W_bits-1 downto 0);

	signal three_xyn_2		: unsigned(W_bits-1 downto 0);

	signal yn_3_xyn_2		: unsigned(2*W_bits-1 downto 0);
	signal yn_3_xyn_2_resized	: unsigned(W_bits-1 downto 0);
	signal yn_3_xyn_2_resized_shift	: unsigned(W_bits-1 downto 0);

	--signal x_test	: std_logic_vector(W_bits-1 downto 0);
	--signal y_test	: std_logic_vector(W_bits-1 downto 0);

	signal delay1	: std_logic_Vector(W_bits-1 downto 0);
	signal delay2	: std_logic_Vector(W_bits-1 downto 0);
	signal delay3	: std_logic_Vector(W_bits-1 downto 0);
	signal delay4	: std_logic_Vector(W_bits-1 downto 0);
	signal delay5	: std_logic_vector(W_bits-1 downto 0);
	signal delay6	: std_logic_vector(W_bits-1 downto 0);
	signal delay7	: std_logic_vector(W_bits-1 downto 0);
	signal delay8	: std_logic_vector(W_bits-1 downto 0);
	signal delay9	: std_logic_vector(W_bits-1 downto 0);
	signal delay10	: std_logic_vector(W_bits-1 downto 0);
	signal delay11	: std_logic_vector(W_bits-1 downto 0);
	signal delay12	: std_logic_vector(W_bits-1 downto 0);

	begin
	


	process(clock)

	begin

	three <= "00000000000000110000000000000000";

	if(rising_edge(clock)) then
	--		yn^2			--

	yn_squared <= unsigned(y_0) * unsigned(y_0);
	
	yn_squared_resized <= yn_squared(W_bits-1+F_bits downto F_bits);

	------------------------------------------

	--		x*yn^2			--

	delay1 <= x;
	delay2 <= delay1;
	delay3 <= delay2;
	delay4 <= delay3;
	delay5 <= delay4;
	delay6 <= delay5;
	delay7 <= delay6;
	delay8 <= delay7;
	delay9 <= delay8;
	delay10<= delay9;
	delay11<= delay10;

	x_test <= delay11;
	

	x_yn_2 <= yn_squared_resized * unsigned(delay11);

	x_yn_2_resized <= x_yn_2(W_bits-1+F_bits downto F_bits);

	------------------------------------------

	--		3-x*yn^2		--

	three_xyn_2 <= unsigned(three) - x_yn_2_resized;


	------------------------------------------
	
	--		yn(3-x*yn^2)		--

	y_test <= y_0;
	yn_3_xyn_2 <= unsigned(y_0)*three_xyn_2;

	yn_3_xyn_2_resized <= yn_3_xyn_2(W_bits-1+F_bits downto F_bits);
	

	------------------------------------------

	--		(yn(3-x*yn*2))/2	--

	yn_3_xyn_2_resized_shift <= shift_right(yn_3_xyn_2_resized,1);

	------------------------------------------


	y <= std_logic_vector(yn_3_xyn_2_resized_shift);
	end if;	
	end process;
end architecture;

