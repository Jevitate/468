
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_unsigned.all;


entity alpha_computation is 
	
	generic(
		W_bits			: positive := 32; -- size of word
		F_bits			: positive := 16); -- number of newton's iterations
		
	port(	clock		: in std_logic;
		beta		: in unsigned(W_bits-1 downto 0);
		alpha		: out unsigned(W_bits-1 downto 0));
		
end entity alpha_computation;



architecture alpha_comp_arch of alpha_computation is

	---- Beta Even, Alpha = -2B + .5B + .5    -- Beta Even Alpha = -2*B + .5*B


	signal beta_one		: unsigned(W_bits-1 downto 0);
	signal beta_two		: unsigned(W_bits-1 downto 0);

	signal even_odd		: std_logic := '0';

	begin
	

	process(clock)

	begin

		if(rising_edge(clock)) then
			if(beta(0) = '1') then -- '1' is odd, '0' is even
				even_odd <= '1';
			elsif(beta(0) = '0') then
				even_odd <= '0';
			end if;		
		
		end if;

	end process;
	
	process(even_odd,clock)

	begin
	if(rising_edge(clock)) then

	beta_one <= shift_left(beta,1);
	beta_two <= shift_right(beta,1);
		if(even_odd = '0') then -- EVEN	
			alpha <= beta_two - beta_one;
		else			 -- ODD
			alpha <= beta_two - beta_one + 1;
		end if;
	end if;
	end process;
	
end architecture;